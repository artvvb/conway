`timescale 1ns / 1ps
module memory_control_sim;
endmodule