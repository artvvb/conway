`timescale 1ns / 1ps
`include "hdl/memory_control.v"
module memory_control_tb;
    wire a;
endmodule