`timescale 1ns / 1ps
`default_nettype none

module data_path (
    input wire clk,
    input wire resetn
);
    
endmodule