`timescale 1ns / 1ps
`include "hdl/data_path.v"
module data_path_tb;
endmodule