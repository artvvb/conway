`timescale 1ns / 1ps
module data_path_sim;
endmodule